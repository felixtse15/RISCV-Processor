module piperegD_Ex(input  logic 	   clk, reset,
				   input  logic 	   clear,
				   input  logic [4:0]  Rs1D, Rs2D, RdD,
				   input  logic [31:0] RD1D, RD2D, PCD, PCPlus4D,
				   input  logic [31:0] ImmExtD,
				   output logic [4:0]  Rs1E, Rs2E, RdE,
				   output logic [31:0] RD1E, RD2E, PCE, PCPlus4E,
				   output logic [31:0] ImmExtE);

	always_ff @ (posedge clk or posedge reset) begin
		if (reset) begin
			RD1E 	 <= 0;
			RD2E 	 <= 0;
			Rs1E 	 <= 0;
			Rs2E     <= 0;
			RdE      <= 0;
			PCE      <= 0;
			PCPlus4E <= 0;
			ImmExtE  <= 0;
		end
		else if (clear) begin
			RD1E 	 <= 0;
			RD2E 	 <= 0;
			Rs1E 	 <= 0;
			Rs2E     <= 0;
			RdE      <= 0;
			PCE      <= 0;
			PCPlus4E <= 0;
			ImmExtE  <= 0;
		end
		else begin
			RD1E 	 <= RD1D;
			RD2E 	 <= RD2D;
			Rs1E 	 <= Rs1D;
			Rs2E     <= Rs2D;
			RdE      <= RdD;
			PCE      <= PCD;
			PCPlus4E <= PCPlus4D;
			ImmExtE  <= ImmExtD;
		end
	end	
	
endmodule